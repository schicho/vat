module printer

const buf_size = 64 * 1024

interface Printer {
	print()
}
